# ====================================================================
#
#      hal_riscv_riscv32.cdl
#
#      RISCV 32 variant architectural HAL package configuration data
#
# ====================================================================
## ####ECOSGPLCOPYRIGHTBEGIN####                                            
## -------------------------------------------                              
## This file is part of eCos, the Embedded Configurable Operating System.   
## Copyright (C) 1998, 1999, 2000, 2001, 2002 Free Software Foundation, Inc.
##
## eCos is free software; you can redistribute it and/or modify it under    
## the terms of the GNU General Public License as published by the Free     
## Software Foundation; either version 2 or (at your option) any later      
## version.                                                                 
##
## eCos is distributed in the hope that it will be useful, but WITHOUT      
## ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or    
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License    
## for more details.                                                        
##
## You should have received a copy of the GNU General Public License        
## along with eCos; if not, write to the Free Software Foundation, Inc.,    
## 51 Franklin Street, Fifth Floor, Boston, MA  02110-1301, USA.            
##
## As a special exception, if other files instantiate templates or use      
## macros or inline functions from this file, or you compile this file      
## and link it with other works to produce a work based on this file,       
## this file does not by itself cause the resulting work to be covered by   
## the GNU General Public License. However the source code for this file    
## must still be made available in accordance with section (3) of the GNU   
## General Public License v2.                                               
##
## This exception does not invalidate any other reasons why a work based    
## on this file might be covered by the GNU General Public License.         
## -------------------------------------------                              
## ####ECOSGPLCOPYRIGHTEND####                                              
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      grihey
# Original data:  grihey
# Contributors:
# Date:           2017-03-17
#
#####DESCRIPTIONEND####
#
# ====================================================================

cdl_package CYGPKG_HAL_RISCV_RISCV32 {
    display       "RISCV32 variant"
    parent        CYGPKG_HAL_RISCV
    hardware
    include_dir   cyg/hal
    description   "
           The RISCV32 architecture HAL package provides generic support
           for this processor architecture. It is also necessary to
           select a specific target platform HAL package."

    cdl_option CYGHWR_HAL_RISCV_RISCV32_CORE {
        display       "RISCV32 processor core used"
        flavor        data
        default_value {"SCR5"}
        legal_values  {"SCR5"}
        description   "
            The RISCV 32 cores." 
    }

    implements    CYGINT_HAL_RISCV_VARIANT

    cdl_option CYGHWR_HAL_RISCV_FPU {
        display    "Variant FPU support"
        calculated 0
    }
    
    cdl_option  CYGHWR_HAL_RISCV_CPU_FREQ {
        display "Variant frequency"
        flavor data
        default_value {"20000000"}
        define -file system.h CYGHWR_HAL_RISCV_CPU_FREQ 
    }
    
    define_proc {
        puts $::cdl_header "#include <pkgconf/hal_riscv.h>"
    }

    compile       var_misc.c variant.S

    make {
        <PREFIX>/lib/target.ld: <PACKAGE>/src/riscv_riscv32.ld
        $(CC) -E -P -Wp,-MD,target.tmp -DEXTRAS=1 -xc $(INCLUDE_PATH) $(CFLAGS) -o $@ $<
        @echo $@ ": \\" > $(notdir $@).deps
        @tail -n +2 target.tmp >> $(notdir $@).deps
        @echo >> $(notdir $@).deps
        @rm target.tmp
    }

    cdl_option CYGBLD_LINKER_SCRIPT {
        display "Linker script"
        flavor data
	no_define
        calculated  { "src/riscv_riscv32.ld" }
    }


    cdl_component CYGBLD_GLOBAL_OPTIONS {
        display "Global build options"
        flavor  none
        parent  CYGPKG_NONE
        description   "
	    Global build options including control over
	    compiler flags, linker flags and choice of toolchain."


        cdl_option CYGBLD_GLOBAL_COMMAND_PREFIX {
            display "Global command prefix"
            flavor  data
            no_define
            default_value { "riscv32-unknown-elf" }
            description "
                This option specifies the command prefix used when
                invoking the build tools."
        }

        cdl_option CYGBLD_GLOBAL_CFLAGS {
            display "Global compiler flags"
            flavor  data
            no_define

            # TODO: add march FPU parameterizing

            default_value { CYGBLD_GLOBAL_WARNFLAGS .
                            "-march=RV32IMA -m32 -std=gnu99 -O2 " .                                                
                            "-fomit-frame-pointer -fno-exceptions -fno-asynchronous-unwind-tables " .
                            "-fno-unwind-tables -fdata-sections -ffunction-sections -fno-common -fno-builtin-printf"
            }
            description   "
                This option controls the global compiler flags which
                are used to compile all packages by
                default. Individual packages may define
                options which override these global flags."
        }

        cdl_option CYGBLD_GLOBAL_LDFLAGS {
            display "Global linker flags"
            flavor  data
            no_define
            default_value { "-static -nostdlib -nostartfiles -Wl,--gc-sections" }
            description   "
                This option controls the global linker flags. Individual
                packages may define options which override these global flags."
        }
    }
}
