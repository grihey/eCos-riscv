# ====================================================================
#
#      hal_riscv_bemicrocva9.cdl
#
#      RISCV BeMicroCV-A9 board HAL package configuration data
#
# ====================================================================
## ####ECOSGPLCOPYRIGHTBEGIN####                                            
## -------------------------------------------                              
## This file is part of eCos, the Embedded Configurable Operating System.   
## Copyright (C) 1998, 1999, 2000, 2001, 2002 Free Software Foundation, Inc.
##
## eCos is free software; you can redistribute it and/or modify it under    
## the terms of the GNU General Public License as published by the Free     
## Software Foundation; either version 2 or (at your option) any later      
## version.                                                                 
##
## eCos is distributed in the hope that it will be useful, but WITHOUT      
## ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or    
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License    
## for more details.                                                        
##
## You should have received a copy of the GNU General Public License        
## along with eCos; if not, write to the Free Software Foundation, Inc.,    
## 51 Franklin Street, Fifth Floor, Boston, MA  02110-1301, USA.            
##
## As a special exception, if other files instantiate templates or use      
## macros or inline functions from this file, or you compile this file      
## and link it with other works to produce a work based on this file,       
## this file does not by itself cause the resulting work to be covered by   
## the GNU General Public License. However the source code for this file    
## must still be made available in accordance with section (3) of the GNU   
## General Public License v2.                                               
##
## This exception does not invalidate any other reasons why a work based    
## on this file might be covered by the GNU General Public License.         
## -------------------------------------------                              
## ####ECOSGPLCOPYRIGHTEND####                                              
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      grihey
# Original data:  bartv
# Contributors:   grihey
# Date:           2017-03-17
#
#####DESCRIPTIONEND####
#
# ====================================================================

cdl_package CYGPKG_HAL_RISCV_BEMICROCVA9 {
    display  "BeMicroCV-A9 board"
    parent        CYGPKG_HAL_RISCV
    define_header   bemicrocva9.h
    include_dir     cyg/hal
    requires      { 
                       (CYGHWR_HAL_RISCV_RISCV32_CORE == "SCR5") && CYGPKG_HAL_RISCV_RISCV32
                  }
    description   "
           The BeMicroCV-A9 HAL package should be used when targetting the
           actual hardware."

    compile       platform.S plf_misc.c hal_diag.c

    cdl_option CYGBLD_HAL_TARGET_H {
        display       "Variant header"
        flavor        data
	    no_define

	calculated { CYGPKG_HAL_RISCV_RISCV32 ? "<pkgconf/hal_riscv_riscv32.h>" : \
                                              "<pkgconf/hal_riscv_riscv64.h>" }
	define -file system.h CYGBLD_HAL_TARGET_H
        description   "Variant header."

        define_proc {
            puts $::cdl_system_header "#define CYGBLD_HAL_PLATFORM_H <pkgconf/bemicrocva9.h>"
            puts $::cdl_system_header ""
            puts $::cdl_system_header "/* Make sure we get the CORE type definitions for HAL_PLATFORM_CPU */"
            puts $::cdl_system_header "#include CYGBLD_HAL_TARGET_H"
            puts $::cdl_system_header "#include CYGBLD_HAL_PLATFORM_H"
	    puts $::cdl_system_header "#define HAL_PLATFORM_BOARD    \"BeMicroCV-A9\""
	    puts $::cdl_system_header "#define HAL_PLATFORM_EXTRA    \"\""
	    puts $::cdl_system_header ""
        puts $::cdl_system_header "#if defined(CYGHWR_HAL_RISCV_RISCV32_CORE_SCR5)"
	    puts $::cdl_system_header "#  define HAL_PLATFORM_CPU    \"RISCV32 SCR5\""
	    puts $::cdl_system_header "#else"
	    puts $::cdl_system_header "#  error Unknown Core"
	    puts $::cdl_system_header "#endif"
	    puts $::cdl_system_header ""
        }
				      
    }

    cdl_component CYG_HAL_STARTUP {
        display       "Startup type"
        flavor        data
        legal_values  {"RAM" "ROM"}
        default_value {"RAM"}
	    no_define
	    define -file system.h CYG_HAL_STARTUP
        description   "
            Currently only ROM startup type is supported."
    }

    cdl_component CYGHWR_UART0_SETTINGS {
        display "uart0 settings"
        no_define
        flavor none
        
        cdl_option CYGHWR_UART0_BASE {
            display         "uart0 base address"
            flavor          data
            default_value   {"0x7fff1200"}
            define CYGHWR_UART0_BASE
        }

        cdl_option CYGHWR_UART0_BAUDRATE {
            display         "uart0 baudrate"
            flavor          data
            default_value   {"115200"}
            define CYGHWR_UART0_BAUDRATE
        }

        cdl_option CYGHWR_UART0_TYPE {
            display         "uart0 controller type"
            flavor          data
            default_value   {"16550"}
            legal_values    {"16450" "16550"}
            define CYGHWR_UART0_TYPE
        }
    }

    # The "-o file" is a workaround for CR100958 - without it the
    # output file would end up in the source directory under CygWin.
    # n.b. grep does not behave itself under win32
    make -priority 1 {
        <PREFIX>/include/cyg/hal/plf_defs.inc : <PACKAGE>/src/plf_mk_defs.c
        $(CC) -E -P -Wp,-MD,target.tmp -DEXTRAS=1 -xc $(INCLUDE_PATH) $(CFLAGS) -o $@ $<
        fgrep .equ plf_mk_defs.tmp | sed s/#// > $@
        @echo $@ ": \\" > $(notdir $@).deps
        @tail -n +2 plf_defs.tmp >> $(notdir $@).deps
        @echo >> $(notdir $@).deps
        @rm plf_defs.tmp plf_mk_defs.tmp
    }

    cdl_option CYGNUM_HAL_VIRTUAL_VECTOR_COMM_CHANNELS {
        display      "Number of communication channels on the board"
        flavor       data
        calculated   1
    }

    cdl_option CYGNUM_HAL_VIRTUAL_VECTOR_DEBUG_CHANNEL {
        display          "Debug serial port"
        active_if        CYGPRI_HAL_VIRTUAL_VECTOR_DEBUG_CHANNEL_CONFIGURABLE
        flavor data
        legal_values     0 to CYGNUM_HAL_VIRTUAL_VECTOR_COMM_CHANNELS-1
        default_value    0
        description      "
           ."
    }

    cdl_option  CYGHWR_HAL_RISCV_CPU_FREQ {
        display "Variant frequency"
        flavor data
        default_value {"20000000"}
        define -file system.h CYGHWR_HAL_RISCV_CPU_FREQ 
    }

    cdl_component CYGNUM_HAL_RTC_CONSTANTS {
        display       "Real-time clock constants."
        flavor        none
    
        cdl_option CYGNUM_HAL_RTC_NUMERATOR {
            display       "Real-time clock numerator"
            flavor        data
            default_value 1000000000
        }
        cdl_option CYGNUM_HAL_RTC_DENOMINATOR {
            display       "Real-time clock denominator"
            flavor        data
            default_value 100
        }
        cdl_option CYGNUM_HAL_RTC_PERIOD {
            display       "Real-time clock period"
            flavor        data
            default_value { ( CYGHWR_HAL_RISCV_CPU_FREQ / 2) / CYGNUM_HAL_RTC_DENOMINATOR }
            description   "
                The count and compare registers of the bemicrocva9 are used
                to drive the eCos kernel RTC. The count register
                increments at half the CPU clock speed."
        }
    }

    cdl_component CYGHWR_MEMORY_LAYOUT {
        display "Memory layout"
        flavor data
        no_define
        calculated { CYG_HAL_STARTUP == "RAM" ? "riscv_bemicrocva9_ram" : \
                                                "riscv_bemicrocva9_rom" }

        cdl_option CYGHWR_MEMORY_LAYOUT_LDI {
            display "Memory layout linker script fragment"
            flavor data
            no_define
            define -file system.h CYGHWR_MEMORY_LAYOUT_LDI
            calculated { CYG_HAL_STARTUP == "RAM" ? "<pkgconf/mlt_riscv_bemicrocva9_ram.ldi>" : \
                                                    "<pkgconf/mlt_riscv_bemicrocva9_rom.ldi>" }
        }

        cdl_option CYGHWR_MEMORY_LAYOUT_H {
            display "Memory layout header file"
            flavor data
            no_define
            define -file system.h CYGHWR_MEMORY_LAYOUT_H
            calculated { CYG_HAL_STARTUP == "RAM" ? "<pkgconf/mlt_riscv_bemicrocva9_ram.h>" : \
                                                    "<pkgconf/mlt_riscv_bemicrocva9_rom.h>" }
        }
    }
}
